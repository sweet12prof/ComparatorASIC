----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    05:21:01 03/27/2020 
-- Design Name: 
-- Module Name:    GreaterComparator - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity GreaterComparator is
	port(
			A,B : in std_logic_vector(7 downto 0);
			greater : out std_logic
		);
end GreaterComparator;

architecture Behavioral of GreaterComparator is

begin
	greater <= '1' when (A > B) else '0';
end Behavioral;

